module subtractor(
	input 		i_a,
	input		i_b,
	output reg	o_y
	);

	assign o_y = i_a - i_b; 

endmodule
