module NOT_gate(
	i_a,
	o_y
	);
	assign o_y = !i_a;
endmodule
